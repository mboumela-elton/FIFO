LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE work.my_package.ALL;

CONFIGURATION cfg_sequenceur OF sequenceur IS
    FOR 